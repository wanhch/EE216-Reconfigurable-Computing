module FIR (
    input  [7:0] din,
    input  clk,
    input  rst,
    output signed [16:0] dout);

    parameter signed [4:0] h0 = 5'd1;
    parameter signed [4:0] h1 = -5'd2;
    parameter signed [4:0] h2 = 5'd3;
    parameter signed [4:0] h3 = -5'd4;
    parameter signed [4:0] h4 = 5'd5;
    parameter signed [4:0] h5 = -5'd6;
    parameter signed [4:0] h6 = 5'd7;
    parameter signed [4:0] h7 = -5'd8;

    reg [7:0] tmp1;
    reg [7:0] tmp2;
    reg [7:0] tmp3;
    reg [7:0] tmp4;
    reg [7:0] tmp5;
    reg [7:0] tmp6;
    reg [7:0] tmp7;
    reg [7:0] tmp8;
    reg [7:0] tmp9;
    reg [7:0] tmp10;
    reg [7:0] tmp11;
    reg [7:0] tmp12;
    reg [7:0] tmp13;
    reg [7:0] tmp14;
    reg [7:0] tmp15;
    reg [15:0] buffer_1_1;
    reg [15:0] buffer_2_1;
    reg [15:0] buffer_2_2;
    reg [15:0] buffer_3_1;
    reg [15:0] buffer_3_2;
    reg [15:0] buffer_3_3;
    reg [15:0] buffer_4_1;
    reg [15:0] buffer_4_2;
    reg [15:0] buffer_4_3;
    reg [15:0] buffer_4_4;
    reg [15:0] buffer_5_1;
    reg [15:0] buffer_5_2;
    reg [15:0] buffer_5_3;
    reg [15:0] buffer_5_4;
    reg [15:0] buffer_5_5;
    reg [15:0] buffer_6_1;
    reg [15:0] buffer_6_2;
    reg [15:0] buffer_6_3;
    reg [15:0] buffer_6_4;
    reg [15:0] buffer_6_5;
    reg [15:0] buffer_6_6;
    reg [15:0] buffer_7_1;
    reg [15:0] buffer_7_2;
    reg [15:0] buffer_7_3;
    reg [15:0] buffer_7_4;
    reg [15:0] buffer_7_5;
    reg [15:0] buffer_7_6;
    reg [15:0] buffer_7_7;
    reg [15:0] buffer_8_1;
    reg [15:0] buffer_8_2;
    reg [15:0] buffer_8_3;
    reg [15:0] buffer_8_4;
    reg [15:0] buffer_8_5;
    reg [15:0] buffer_8_6;
    reg [15:0] buffer_8_7;
    reg [15:0] buffer_8_8;
    reg [15:0] buffer_2to3;
    reg [15:0] buffer_3to4;
    reg [15:0] buffer_4to5;
    reg [15:0] buffer_5to6;
    reg [15:0] buffer_6to7;
    reg [15:0] buffer_7to8;

    wire [7:0] input1_sig;
    wire [7:0] input2_sig;
    wire [7:0] input3_sig;
    wire [7:0] input4_sig;
    wire [7:0] input5_sig;
    wire [7:0] input6_sig;
    wire [7:0] input7_sig;
    wire [7:0] input8_sig;
    wire [7:0] input9_sig;
    wire [7:0] input10_sig;
    wire [7:0] input11_sig;
    wire [7:0] input12_sig;
    wire [7:0] input13_sig;
    wire [7:0] input14_sig;
    wire [7:0] input15_sig;
    wire [7:0] input16_sig;
    wire [15:0] A1_sig;
    wire [15:0] A2_sig;
    wire [15:0] A3_sig;
    wire [15:0] A4_sig;
    wire [15:0] A5_sig;
    wire [15:0] A6_sig;
    wire [15:0] A7_sig;
    wire [15:0] A8_sig;
    wire [15:0] M1_sig;
    wire [15:0] M2_sig;
    wire [15:0] M3_sig;
    wire [15:0] M4_sig;
    wire [15:0] M5_sig;
    wire [15:0] M6_sig;
    wire [15:0] M7_sig;
    wire [15:0] M8_sig;

    wire [15:0] buffered_M1_sig;
    wire [15:0] buffered_M2_sig;
    wire [15:0] buffered_M3_sig;
    wire [15:0] buffered_M4_sig;
    wire [15:0] buffered_M5_sig;
    wire [15:0] buffered_M6_sig;
    wire [15:0] buffered_M7_sig;
    wire [15:0] buffered_M8_sig;

    wire [15:0] CA_2_sig;
    wire [15:0] CA_3_sig;
    wire [15:0] CA_4_sig;
    wire [15:0] CA_5_sig;
    wire [15:0] CA_6_sig;
    wire [15:0] CA_7_sig;
    wire [15:0] CA_2_buffered_sig;
    wire [15:0] CA_3_buffered_sig;
    wire [15:0] CA_4_buffered_sig;
    wire [15:0] CA_5_buffered_sig;
    wire [15:0] CA_6_buffered_sig;
    wire [15:0] CA_7_buffered_sig;

    assign input1_sig = din;
    assign input2_sig = tmp1;
    assign input3_sig = tmp2;
    assign input4_sig = tmp3;
    assign input5_sig = tmp4;
    assign input6_sig = tmp5;
    assign input7_sig = tmp6;
    assign input8_sig = tmp7;
    assign input9_sig = tmp8;
    assign input10_sig = tmp9;
    assign input11_sig = tmp10;
    assign input12_sig = tmp11;
    assign input13_sig = tmp12;
    assign input14_sig = tmp13;
    assign input15_sig = tmp14;
    assign input16_sig = tmp15;

    MultiCycleAdder MA_1(input1_sig, input16_sig, 0, clk, rst, A1_sig);
    MultiCycleAdder MA_2(input2_sig, input15_sig, 0, clk, rst, A2_sig);
    MultiCycleAdder MA_3(input3_sig, input14_sig, 0, clk, rst, A3_sig);
    MultiCycleAdder MA_4(input4_sig, input13_sig, 0, clk, rst, A4_sig);
    MultiCycleAdder MA_5(input5_sig, input12_sig, 0, clk, rst, A5_sig);
    MultiCycleAdder MA_6(input6_sig, input11_sig, 0, clk, rst, A6_sig);
    MultiCycleAdder MA_7(input7_sig, input10_sig, 0, clk, rst, A7_sig);
    MultiCycleAdder MA_8(input8_sig, input9_sig, 0, clk, rst, A8_sig);

    assign buffered_M1_sig = buffer_1_1;
    assign buffered_M2_sig = buffer_2_1;
    assign buffered_M3_sig = buffer_3_2;
    assign buffered_M4_sig = buffer_4_3;
    assign buffered_M5_sig = buffer_5_4;
    assign buffered_M6_sig = buffer_6_5;
    assign buffered_M7_sig = buffer_7_6;
    assign buffered_M8_sig = buffer_8_7;

    assign CA_2_buffered_sig = buffer_2to3;
    assign CA_3_buffered_sig = buffer_3to4;
    assign CA_4_buffered_sig = buffer_4to5;
    assign CA_5_buffered_sig = buffer_5to6;
    assign CA_6_buffered_sig = buffer_6to7;
    assign CA_7_buffered_sig = buffer_7to8;

    MultiCycleAdder CA_2(buffered_M1_sig, buffered_M2_sig, 0, clk, rst, CA_2_sig);
    MultiCycleAdder CA_3(CA_2_buffered_sig, buffered_M3_sig, 0, clk, rst, CA_3_sig);
    MultiCycleAdder CA_4(CA_3_buffered_sig, buffered_M4_sig, 0, clk, rst, CA_4_sig);
    MultiCycleAdder CA_5(CA_4_buffered_sig, buffered_M5_sig, 0, clk, rst, CA_5_sig);
    MultiCycleAdder CA_6(CA_5_buffered_sig, buffered_M6_sig, 0, clk, rst, CA_6_sig);
    MultiCycleAdder CA_7(CA_6_buffered_sig, buffered_M7_sig, 0, clk, rst, CA_7_sig);
    MultiCycleAdder CA_8(CA_7_buffered_sig, buffered_M8_sig, 0, clk, rst, dout);

    always @(posedge clk, posedge rst) begin
        if (rst == 1'b0) begin
            tmp1 <= 8'd0;
            tmp2 <= 8'd0;
            tmp3 <= 8'd0;
            tmp4 <= 8'd0;
            tmp5 <= 8'd0;
            tmp6 <= 8'd0;
            tmp7 <= 8'd0;
            tmp8 <= 8'd0;
            tmp9 <= 8'd0;
            tmp10 <= 8'd0;
            tmp11 <= 8'd0;
            tmp12 <= 8'd0;
            tmp13 <= 8'd0;
            tmp14 <= 8'd0;
            tmp15 <= 8'd0;

            buffer_1_1 <= 16'd0;
            buffer_2_1 <= 16'd0;
            buffer_3_1 <= 16'd0;
            buffer_4_1 <= 16'd0;
            buffer_5_1 <= 16'd0;
            buffer_6_1 <= 16'd0;
            buffer_7_1 <= 16'd0;
            buffer_8_1 <= 16'd0;
            buffer_2_2 <= 16'd0;
            buffer_3_2 <= 16'd0;
            buffer_4_2 <= 16'd0;
            buffer_5_2 <= 16'd0;
            buffer_6_2 <= 16'd0;
            buffer_7_2 <= 16'd0;
            buffer_8_2 <= 16'd0;
            buffer_3_3 <= 16'd0;
            buffer_4_3 <= 16'd0;
            buffer_5_3 <= 16'd0;
            buffer_6_3 <= 16'd0;
            buffer_7_3 <= 16'd0;
            buffer_8_3 <= 16'd0;
            buffer_4_4 <= 16'd0;
            buffer_5_4 <= 16'd0;
            buffer_6_4 <= 16'd0;
            buffer_7_4 <= 16'd0;
            buffer_8_4 <= 16'd0;
            buffer_5_5 <= 16'd0;
            buffer_6_5 <= 16'd0;
            buffer_7_5 <= 16'd0;
            buffer_8_5 <= 16'd0;
            buffer_6_6 <= 16'd0;
            buffer_7_6 <= 16'd0;
            buffer_8_6 <= 16'd0;
            buffer_7_7 <= 16'd0;
            buffer_8_7 <= 16'd0;
            buffer_8_8 <= 16'd0;

            buffer_2to3 <= 16'd0;
            buffer_3to4 <= 16'd0;
            buffer_4to5 <= 16'd0;
            buffer_5to6 <= 16'd0;
            buffer_6to7 <= 16'd0;
            buffer_7to8 <= 16'd0;
        end else begin
            tmp1 <= din;
            tmp2 <= tmp1;
            tmp3 <= tmp2;
            tmp4 <= tmp3;
            tmp5 <= tmp4;
            tmp6 <= tmp5;
            tmp7 <= tmp6;
            tmp8 <= tmp7;
            tmp9 <= tmp8;
            tmp10 <= tmp9;
            tmp11 <= tmp10;
            tmp12 <= tmp11;
            tmp13 <= tmp12;
            tmp14 <= tmp13;
            tmp15 <= tmp14;

            buffer_1_1 <= A1_sig * h0;
            buffer_2_1 <= A2_sig * h1;
            buffer_3_1 <= A3_sig * h2;
            buffer_4_1 <= A4_sig * h3;
            buffer_5_1 <= A5_sig * h4;
            buffer_6_1 <= A6_sig * h5;
            buffer_7_1 <= A7_sig * h6;
            buffer_8_1 <= A8_sig * h7;
            buffer_2_2 <= buffer_2_1;
            buffer_3_2 <= buffer_3_1;
            buffer_4_2 <= buffer_4_1;
            buffer_5_2 <= buffer_5_1;
            buffer_6_2 <= buffer_6_1;
            buffer_7_2 <= buffer_7_1;
            buffer_8_2 <= buffer_8_1;
            buffer_3_3 <= buffer_3_2;
            buffer_4_3 <= buffer_4_2;
            buffer_5_3 <= buffer_5_2;
            buffer_6_3 <= buffer_6_2;
            buffer_7_3 <= buffer_7_2;
            buffer_8_3 <= buffer_8_2;
            buffer_4_4 <= buffer_4_3;
            buffer_5_4 <= buffer_5_3;
            buffer_6_4 <= buffer_6_3;
            buffer_7_4 <= buffer_7_3;
            buffer_8_4 <= buffer_8_3;
            buffer_5_5 <= buffer_5_4;
            buffer_6_5 <= buffer_6_4;
            buffer_7_5 <= buffer_7_4;
            buffer_8_5 <= buffer_8_4;
            buffer_6_6 <= buffer_6_5;
            buffer_7_6 <= buffer_7_5;
            buffer_8_6 <= buffer_8_5;
            buffer_7_7 <= buffer_7_6;
            buffer_8_7 <= buffer_8_6;
            buffer_8_8 <= buffer_8_7;

            buffer_2to3 <= CA_2_sig;
            buffer_3to4 <= CA_3_sig;
            buffer_4to5 <= CA_4_sig;
            buffer_5to6 <= CA_5_sig;
            buffer_6to7 <= CA_6_sig;
            buffer_7to8 <= CA_7_sig;
        end
    end
endmodule